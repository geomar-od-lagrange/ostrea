netcdf \15m_ds_conn_14 {
dimensions:
	hex0 = 8223 ;
	hex1 = 8282 ;
	month = 5 ;
	year = 4 ;
	corner = 7 ;
variables:
	double aqc_count_hex0(hex0) ;
		aqc_count_hex0:_FillValue = NaN ;
		aqc_count_hex0:coordinates = "hex_label lat_hex0 lon_hex0" ;
	double rst_count_hex0(hex0) ;
		rst_count_hex0:_FillValue = NaN ;
		rst_count_hex0:coordinates = "hex_label lat_hex0 lon_hex0" ;
	double pop_count_hex0(hex0) ;
		pop_count_hex0:_FillValue = NaN ;
		pop_count_hex0:coordinates = "hex_label lat_hex0 lon_hex0" ;
	double dss_count_hex0(hex0) ;
		dss_count_hex0:_FillValue = NaN ;
		dss_count_hex0:coordinates = "hex_label lat_hex0 lon_hex0" ;
	double hly_count_hex0(hex0) ;
		hly_count_hex0:_FillValue = NaN ;
		hly_count_hex0:coordinates = "hex_label lat_hex0 lon_hex0" ;
	double his_count_hex0(hex0) ;
		his_count_hex0:_FillValue = NaN ;
		his_count_hex0:coordinates = "hex_label lat_hex0 lon_hex0" ;
	double aqc_count_hex1(hex1) ;
		aqc_count_hex1:_FillValue = NaN ;
		aqc_count_hex1:coordinates = "lat_hex1 lon_hex1" ;
	double rst_count_hex1(hex1) ;
		rst_count_hex1:_FillValue = NaN ;
		rst_count_hex1:coordinates = "lat_hex1 lon_hex1" ;
	double pop_count_hex1(hex1) ;
		pop_count_hex1:_FillValue = NaN ;
		pop_count_hex1:coordinates = "lat_hex1 lon_hex1" ;
	double dss_count_hex1(hex1) ;
		dss_count_hex1:_FillValue = NaN ;
		dss_count_hex1:coordinates = "lat_hex1 lon_hex1" ;
	double hly_count_hex1(hex1) ;
		hly_count_hex1:_FillValue = NaN ;
		hly_count_hex1:coordinates = "lat_hex1 lon_hex1" ;
	double his_count_hex1(hex1) ;
		his_count_hex1:_FillValue = NaN ;
		his_count_hex1:coordinates = "lat_hex1 lon_hex1" ;
	double obs(month, year, hex0, hex1) ;
		obs:_FillValue = NaN ;
		obs:coordinates = "hex_label lat_hex0 lat_hex1 lon_hex0 lon_hex1" ;
	double water_fraction_hex0(hex0) ;
		water_fraction_hex0:_FillValue = NaN ;
		water_fraction_hex0:coordinates = "hex_label lat_hex0 lon_hex0" ;
	double water_fraction_hex1(hex1) ;
		water_fraction_hex1:_FillValue = NaN ;
		water_fraction_hex1:coordinates = "lat_hex1 lon_hex1" ;
	float gridbox_count_hex0(hex0) ;
		gridbox_count_hex0:_FillValue = NaNf ;
		gridbox_count_hex0:coordinates = "hex_label lat_hex0 lon_hex0" ;
	float gridbox_count_hex1(hex1) ;
		gridbox_count_hex1:_FillValue = NaNf ;
		gridbox_count_hex1:coordinates = "lat_hex1 lon_hex1" ;
	double water_count_hex0(hex0) ;
		water_count_hex0:_FillValue = NaN ;
		water_count_hex0:coordinates = "hex_label lat_hex0 lon_hex0" ;
	double water_count_hex1(hex1) ;
		water_count_hex1:_FillValue = NaN ;
		water_count_hex1:coordinates = "lat_hex1 lon_hex1" ;
	float depth_mean_hex0(hex0) ;
		depth_mean_hex0:_FillValue = NaNf ;
		depth_mean_hex0:coordinates = "hex_label lat_hex0 lon_hex0" ;
	float depth_mean_hex1(hex1) ;
		depth_mean_hex1:_FillValue = NaNf ;
		depth_mean_hex1:coordinates = "lat_hex1 lon_hex1" ;
	double depth_median_hex0(hex0) ;
		depth_median_hex0:_FillValue = NaN ;
		depth_median_hex0:coordinates = "hex_label lat_hex0 lon_hex0" ;
	double depth_median_hex1(hex1) ;
		depth_median_hex1:_FillValue = NaN ;
		depth_median_hex1:coordinates = "lat_hex1 lon_hex1" ;
	float depth_std_hex0(hex0) ;
		depth_std_hex0:_FillValue = NaNf ;
		depth_std_hex0:coordinates = "hex_label lat_hex0 lon_hex0" ;
	float depth_std_hex1(hex1) ;
		depth_std_hex1:_FillValue = NaNf ;
		depth_std_hex1:coordinates = "lat_hex1 lon_hex1" ;
	string hex0(hex0) ;
	string hex1(hex1) ;
	double month(month) ;
		month:_FillValue = NaN ;
	double year(year) ;
		year:_FillValue = NaN ;
	double lon_hex0_corners(corner, hex0) ;
		lon_hex0_corners:_FillValue = NaN ;
	double lat_hex0_corners(corner, hex0) ;
		lat_hex0_corners:_FillValue = NaN ;
	double lon_hex1_corners(corner, hex1) ;
		lon_hex1_corners:_FillValue = NaN ;
	double lat_hex1_corners(corner, hex1) ;
		lat_hex1_corners:_FillValue = NaN ;
	double lon_hex0(hex0) ;
		lon_hex0:_FillValue = NaN ;
	double lon_hex1(hex1) ;
		lon_hex1:_FillValue = NaN ;
	double lat_hex0(hex0) ;
		lat_hex0:_FillValue = NaN ;
	double lat_hex1(hex1) ;
		lat_hex1:_FillValue = NaN ;
	string hex_label(hex0) ;
	double obs_per_origin_area(month, year, hex0, hex1) ;
		obs_per_origin_area:_FillValue = NaN ;
		obs_per_origin_area:coordinates = "hex_label lat_hex0 lat_hex1 lon_hex0 lon_hex1" ;
	byte habitable_hex0(hex0) ;
		habitable_hex0:coordinates = "hex_label lat_hex0 lon_hex0" ;
		habitable_hex0:dtype = "bool" ;
	byte habitable_hex1(hex1) ;
		habitable_hex1:coordinates = "lat_hex1 lon_hex1" ;
		habitable_hex1:dtype = "bool" ;

// global attributes:
		:coordinates = "lat_hex0_corners lat_hex1_corners lon_hex0_corners lon_hex1_corners" ;
}
